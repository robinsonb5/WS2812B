-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity WS2812B_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end WS2812B_ROM;

architecture arch of WS2812B_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"84808080",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"40000016",
     7 => x"00000000",
     8 => x"8480808c",
     9 => x"f0088480",
    10 => x"808cf408",
    11 => x"8480808c",
    12 => x"f8088480",
    13 => x"80809808",
    14 => x"2d848080",
    15 => x"8cf80c84",
    16 => x"80808cf4",
    17 => x"0c848080",
    18 => x"8cf00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"80808ce0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"8480808c",
    57 => x"f0708480",
    58 => x"8099e427",
    59 => x"8e388071",
    60 => x"70840553",
    61 => x"0c848080",
    62 => x"81e50484",
    63 => x"8080808c",
    64 => x"51848080",
    65 => x"86fc0402",
    66 => x"f8050d73",
    67 => x"52ff8408",
    68 => x"70882a70",
    69 => x"81065151",
    70 => x"5170802e",
    71 => x"f03871ff",
    72 => x"840c7184",
    73 => x"80808cf0",
    74 => x"0c028805",
    75 => x"0d0402f0",
    76 => x"050d7553",
    77 => x"80738480",
    78 => x"8080f52d",
    79 => x"7081ff06",
    80 => x"53535470",
    81 => x"742eb138",
    82 => x"7181ff06",
    83 => x"81145452",
    84 => x"ff840870",
    85 => x"882a7081",
    86 => x"06515151",
    87 => x"70802ef0",
    88 => x"3871ff84",
    89 => x"0c811473",
    90 => x"84808080",
    91 => x"f52d7081",
    92 => x"ff065353",
    93 => x"5470d138",
    94 => x"73848080",
    95 => x"8cf00c02",
    96 => x"90050d04",
    97 => x"02f8050d",
    98 => x"ff840870",
    99 => x"892a7081",
   100 => x"06515252",
   101 => x"70802ef0",
   102 => x"387181ff",
   103 => x"06848080",
   104 => x"8cf00c02",
   105 => x"88050d04",
   106 => x"02c4050d",
   107 => x"0280c005",
   108 => x"8480808d",
   109 => x"d05b5680",
   110 => x"76708405",
   111 => x"5808715e",
   112 => x"5e577c70",
   113 => x"84055e08",
   114 => x"58805b77",
   115 => x"982a7888",
   116 => x"2b595372",
   117 => x"8938765e",
   118 => x"84808085",
   119 => x"e3047b80",
   120 => x"2e81d838",
   121 => x"805c7280",
   122 => x"e42ea138",
   123 => x"7280e426",
   124 => x"8e387280",
   125 => x"e32e80f5",
   126 => x"38848080",
   127 => x"84fb0472",
   128 => x"80f32e80",
   129 => x"d0388480",
   130 => x"8084fb04",
   131 => x"75841771",
   132 => x"087e5c56",
   133 => x"57528755",
   134 => x"739c2a74",
   135 => x"842b5552",
   136 => x"71802e83",
   137 => x"38815989",
   138 => x"72258a38",
   139 => x"b7125284",
   140 => x"808084b8",
   141 => x"04b01252",
   142 => x"78802e89",
   143 => x"38715184",
   144 => x"80808287",
   145 => x"2dff1555",
   146 => x"748025cc",
   147 => x"38805484",
   148 => x"80808594",
   149 => x"04758417",
   150 => x"71087054",
   151 => x"5c575284",
   152 => x"808082ae",
   153 => x"2d7b5484",
   154 => x"80808594",
   155 => x"04758417",
   156 => x"71085557",
   157 => x"52848080",
   158 => x"85cb04a5",
   159 => x"51848080",
   160 => x"82872d72",
   161 => x"51848080",
   162 => x"82872d82",
   163 => x"17578480",
   164 => x"8085d604",
   165 => x"73ff1555",
   166 => x"52807225",
   167 => x"b9387970",
   168 => x"81055b84",
   169 => x"808080f5",
   170 => x"2d705253",
   171 => x"84808082",
   172 => x"872d8117",
   173 => x"57848080",
   174 => x"85940472",
   175 => x"a52e0981",
   176 => x"06893881",
   177 => x"5c848080",
   178 => x"85d60472",
   179 => x"51848080",
   180 => x"82872d81",
   181 => x"1757811b",
   182 => x"5b837b25",
   183 => x"fded3872",
   184 => x"fde0387d",
   185 => x"8480808c",
   186 => x"f00c02bc",
   187 => x"050d0402",
   188 => x"f8050d73",
   189 => x"51bd5280",
   190 => x"710c800b",
   191 => x"81f8120c",
   192 => x"ff128412",
   193 => x"52527180",
   194 => x"25ed3802",
   195 => x"88050d04",
   196 => x"02e8050d",
   197 => x"77841153",
   198 => x"56bb5571",
   199 => x"0881f813",
   200 => x"08057270",
   201 => x"8405540c",
   202 => x"ff155574",
   203 => x"8025ec38",
   204 => x"81557484",
   205 => x"29167070",
   206 => x"70840552",
   207 => x"08701011",
   208 => x"fc140810",
   209 => x"11730810",
   210 => x"1170832c",
   211 => x"74317083",
   212 => x"2b81f818",
   213 => x"70089029",
   214 => x"71083170",
   215 => x"842c7384",
   216 => x"2c05720c",
   217 => x"58585151",
   218 => x"51515481",
   219 => x"18585654",
   220 => x"52bc7525",
   221 => x"ffbc3802",
   222 => x"98050d04",
   223 => x"02ffb805",
   224 => x"0d848080",
   225 => x"8e905184",
   226 => x"808085ef",
   227 => x"2d848080",
   228 => x"92805184",
   229 => x"808085ef",
   230 => x"2d848080",
   231 => x"95f45184",
   232 => x"808085ef",
   233 => x"2db35981",
   234 => x"c2e60b84",
   235 => x"808095f0",
   236 => x"0c78802e",
   237 => x"8a38ff19",
   238 => x"59848080",
   239 => x"89ea0484",
   240 => x"808095f0",
   241 => x"08107084",
   242 => x"808095f0",
   243 => x"0c70962a",
   244 => x"70810651",
   245 => x"53537180",
   246 => x"2e8a3872",
   247 => x"81078480",
   248 => x"8095f00c",
   249 => x"84808095",
   250 => x"f0087095",
   251 => x"2a708106",
   252 => x"51535371",
   253 => x"802e8a38",
   254 => x"72813284",
   255 => x"808095f0",
   256 => x"0c848080",
   257 => x"95f00870",
   258 => x"bf068105",
   259 => x"5454bb73",
   260 => x"258338bb",
   261 => x"53739fff",
   262 => x"ff065297",
   263 => x"ffff7225",
   264 => x"8b387110",
   265 => x"12ffb880",
   266 => x"80115152",
   267 => x"7183ffff",
   268 => x"248d3883",
   269 => x"ffff725b",
   270 => x"41848080",
   271 => x"88d00471",
   272 => x"87ffff24",
   273 => x"933887ff",
   274 => x"ff723141",
   275 => x"83ffff5a",
   276 => x"78428480",
   277 => x"8089b204",
   278 => x"718bffff",
   279 => x"24933878",
   280 => x"4183ffff",
   281 => x"0bf88080",
   282 => x"13435a84",
   283 => x"808089b2",
   284 => x"04718fff",
   285 => x"ff248f38",
   286 => x"788fffff",
   287 => x"73315b41",
   288 => x"84808089",
   289 => x"94047193",
   290 => x"ffff2492",
   291 => x"38f08080",
   292 => x"12795b41",
   293 => x"83ffff42",
   294 => x"84808089",
   295 => x"b2047197",
   296 => x"ffff248e",
   297 => x"3883ffff",
   298 => x"41800b97",
   299 => x"ffff7331",
   300 => x"435a7282",
   301 => x"2b848080",
   302 => x"8e901108",
   303 => x"62058480",
   304 => x"808e9012",
   305 => x"0c848080",
   306 => x"92801108",
   307 => x"1b848080",
   308 => x"9280120c",
   309 => x"84808095",
   310 => x"f4110863",
   311 => x"05848080",
   312 => x"95f4120c",
   313 => x"527381ff",
   314 => x"0659a787",
   315 => x"58ff8408",
   316 => x"ff195952",
   317 => x"778025f5",
   318 => x"38848080",
   319 => x"95f40b84",
   320 => x"05848080",
   321 => x"92800b84",
   322 => x"05848080",
   323 => x"8e900b84",
   324 => x"0581f813",
   325 => x"81f81381",
   326 => x"f8134040",
   327 => x"40404040",
   328 => x"bb587a08",
   329 => x"9f2c7b08",
   330 => x"9f2c7c08",
   331 => x"32707231",
   332 => x"7e089f2c",
   333 => x"7f089f2c",
   334 => x"60083270",
   335 => x"72316208",
   336 => x"9f2c6308",
   337 => x"9f2c6408",
   338 => x"32707231",
   339 => x"66707084",
   340 => x"05520870",
   341 => x"101169fc",
   342 => x"05081011",
   343 => x"73081011",
   344 => x"70832c74",
   345 => x"3170832b",
   346 => x"51515151",
   347 => x"555e5c51",
   348 => x"5c53515a",
   349 => x"53515852",
   350 => x"7180258b",
   351 => x"38767231",
   352 => x"57848080",
   353 => x"8b8a0471",
   354 => x"17577e70",
   355 => x"70840552",
   356 => x"08701011",
   357 => x"61fc0508",
   358 => x"10117308",
   359 => x"10117083",
   360 => x"2c743170",
   361 => x"832b5651",
   362 => x"51515555",
   363 => x"52718025",
   364 => x"8b387572",
   365 => x"31568480",
   366 => x"808bbf04",
   367 => x"7116567f",
   368 => x"70708405",
   369 => x"52087010",
   370 => x"1162fc05",
   371 => x"08101173",
   372 => x"08101170",
   373 => x"832c7431",
   374 => x"70832b56",
   375 => x"51515155",
   376 => x"55527180",
   377 => x"258b3874",
   378 => x"72315584",
   379 => x"80808bf4",
   380 => x"04711555",
   381 => x"74882c70",
   382 => x"81ff0678",
   383 => x"882b87fc",
   384 => x"80800670",
   385 => x"7983fe80",
   386 => x"06077073",
   387 => x"07fc0c51",
   388 => x"54ff1a84",
   389 => x"1e7f8405",
   390 => x"61840563",
   391 => x"84056584",
   392 => x"05678405",
   393 => x"48464442",
   394 => x"405e5a51",
   395 => x"55778025",
   396 => x"fdf03884",
   397 => x"80808e90",
   398 => x"51848080",
   399 => x"86902d84",
   400 => x"80809280",
   401 => x"51848080",
   402 => x"86902d84",
   403 => x"808095f4",
   404 => x"51848080",
   405 => x"86902d84",
   406 => x"808087b1",
   407 => x"04000000",
   408 => x"00ffffff",
   409 => x"ff00ffff",
   410 => x"ffff00ff",
   411 => x"ffffff00",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

