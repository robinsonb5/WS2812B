-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity WS2812B_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end WS2812B_ROM;

architecture arch of WS2812B_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"84808080",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"40000016",
     7 => x"00000000",
     8 => x"8480809a",
     9 => x"cc088480",
    10 => x"809ad008",
    11 => x"8480809a",
    12 => x"d4088480",
    13 => x"80809808",
    14 => x"2d848080",
    15 => x"9ad40c84",
    16 => x"80809ad0",
    17 => x"0c848080",
    18 => x"9acc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"808098fc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"8480809a",
    57 => x"cc708480",
    58 => x"80b8cc27",
    59 => x"8e388071",
    60 => x"70840553",
    61 => x"0c848080",
    62 => x"81e50484",
    63 => x"8080808c",
    64 => x"51848080",
    65 => x"97a90402",
    66 => x"f8050d73",
    67 => x"52ff8408",
    68 => x"70882a70",
    69 => x"81065151",
    70 => x"5170802e",
    71 => x"f03871ff",
    72 => x"840c7184",
    73 => x"80809acc",
    74 => x"0c028805",
    75 => x"0d0402f0",
    76 => x"050d7553",
    77 => x"80738480",
    78 => x"8080f52d",
    79 => x"7081ff06",
    80 => x"53535470",
    81 => x"742eb138",
    82 => x"7181ff06",
    83 => x"81145452",
    84 => x"ff840870",
    85 => x"882a7081",
    86 => x"06515151",
    87 => x"70802ef0",
    88 => x"3871ff84",
    89 => x"0c811473",
    90 => x"84808080",
    91 => x"f52d7081",
    92 => x"ff065353",
    93 => x"5470d138",
    94 => x"73848080",
    95 => x"9acc0c02",
    96 => x"90050d04",
    97 => x"02f8050d",
    98 => x"ff840870",
    99 => x"892a7081",
   100 => x"06515252",
   101 => x"70802ef0",
   102 => x"387181ff",
   103 => x"06848080",
   104 => x"9acc0c02",
   105 => x"88050d04",
   106 => x"02c4050d",
   107 => x"0280c005",
   108 => x"8480809b",
   109 => x"ac5b5680",
   110 => x"76708405",
   111 => x"5808715e",
   112 => x"5e577c70",
   113 => x"84055e08",
   114 => x"58805b77",
   115 => x"982a7888",
   116 => x"2b595372",
   117 => x"8938765e",
   118 => x"84808085",
   119 => x"e3047b80",
   120 => x"2e81d838",
   121 => x"805c7280",
   122 => x"e42ea138",
   123 => x"7280e426",
   124 => x"8e387280",
   125 => x"e32e80f5",
   126 => x"38848080",
   127 => x"84fb0472",
   128 => x"80f32e80",
   129 => x"d0388480",
   130 => x"8084fb04",
   131 => x"75841771",
   132 => x"087e5c56",
   133 => x"57528755",
   134 => x"739c2a74",
   135 => x"842b5552",
   136 => x"71802e83",
   137 => x"38815989",
   138 => x"72258a38",
   139 => x"b7125284",
   140 => x"808084b8",
   141 => x"04b01252",
   142 => x"78802e89",
   143 => x"38715184",
   144 => x"80808287",
   145 => x"2dff1555",
   146 => x"748025cc",
   147 => x"38805484",
   148 => x"80808594",
   149 => x"04758417",
   150 => x"71087054",
   151 => x"5c575284",
   152 => x"808082ae",
   153 => x"2d7b5484",
   154 => x"80808594",
   155 => x"04758417",
   156 => x"71085557",
   157 => x"52848080",
   158 => x"85cb04a5",
   159 => x"51848080",
   160 => x"82872d72",
   161 => x"51848080",
   162 => x"82872d82",
   163 => x"17578480",
   164 => x"8085d604",
   165 => x"73ff1555",
   166 => x"52807225",
   167 => x"b9387970",
   168 => x"81055b84",
   169 => x"808080f5",
   170 => x"2d705253",
   171 => x"84808082",
   172 => x"872d8117",
   173 => x"57848080",
   174 => x"85940472",
   175 => x"a52e0981",
   176 => x"06893881",
   177 => x"5c848080",
   178 => x"85d60472",
   179 => x"51848080",
   180 => x"82872d81",
   181 => x"1757811b",
   182 => x"5b837b25",
   183 => x"fded3872",
   184 => x"fde0387d",
   185 => x"8480809a",
   186 => x"cc0c02bc",
   187 => x"050d0402",
   188 => x"e8050d78",
   189 => x"84115555",
   190 => x"81955689",
   191 => x"cc140888",
   192 => x"2c938c15",
   193 => x"08882c8c",
   194 => x"1608882c",
   195 => x"77080555",
   196 => x"535181ff",
   197 => x"73258438",
   198 => x"81ff5384",
   199 => x"15081151",
   200 => x"81ff7125",
   201 => x"843881ff",
   202 => x"51881508",
   203 => x"125281ff",
   204 => x"72258438",
   205 => x"81ff5272",
   206 => x"902b7188",
   207 => x"2b077073",
   208 => x"07fc0c51",
   209 => x"ff168415",
   210 => x"55567580",
   211 => x"25ffac38",
   212 => x"0298050d",
   213 => x"0402ec05",
   214 => x"0d76788c",
   215 => x"11547153",
   216 => x"84120855",
   217 => x"5654722d",
   218 => x"89cc1552",
   219 => x"73518414",
   220 => x"0853722d",
   221 => x"938c1552",
   222 => x"73518414",
   223 => x"0853722d",
   224 => x"0294050d",
   225 => x"0402f405",
   226 => x"0d757052",
   227 => x"53819752",
   228 => x"800b8c12",
   229 => x"0c800b84",
   230 => x"ec120c80",
   231 => x"0b89cc12",
   232 => x"0c800b8e",
   233 => x"ac120c80",
   234 => x"0b938c12",
   235 => x"0c800b97",
   236 => x"ec120cff",
   237 => x"12841252",
   238 => x"52718025",
   239 => x"d3388073",
   240 => x"0c800b84",
   241 => x"140c800b",
   242 => x"88140c02",
   243 => x"8c050d04",
   244 => x"02e8050d",
   245 => x"77798480",
   246 => x"809bf808",
   247 => x"55575572",
   248 => x"802e8f38",
   249 => x"ff138480",
   250 => x"809bf80c",
   251 => x"84808088",
   252 => x"ce047552",
   253 => x"74519415",
   254 => x"0853722d",
   255 => x"8480809b",
   256 => x"fc081070",
   257 => x"8480809b",
   258 => x"fc0c7096",
   259 => x"2a708106",
   260 => x"51545472",
   261 => x"802e8a38",
   262 => x"73810784",
   263 => x"80809bfc",
   264 => x"0c848080",
   265 => x"9bfc0870",
   266 => x"952a7081",
   267 => x"06515454",
   268 => x"72802e8a",
   269 => x"38738132",
   270 => x"8480809b",
   271 => x"fc0c8480",
   272 => x"809bfc08",
   273 => x"98160806",
   274 => x"8480809b",
   275 => x"f80c7552",
   276 => x"74518815",
   277 => x"0853722d",
   278 => x"0298050d",
   279 => x"0402f005",
   280 => x"0d757779",
   281 => x"7b575553",
   282 => x"5197ffff",
   283 => x"71258b38",
   284 => x"701011ff",
   285 => x"b8808011",
   286 => x"51517083",
   287 => x"ffff248f",
   288 => x"3883ffff",
   289 => x"720c7073",
   290 => x"0c848080",
   291 => x"89a20470",
   292 => x"87ffff24",
   293 => x"963887ff",
   294 => x"ff713172",
   295 => x"0c83ffff",
   296 => x"730c8074",
   297 => x"0c848080",
   298 => x"8a8e0470",
   299 => x"8bffff24",
   300 => x"95388072",
   301 => x"0c83ffff",
   302 => x"730cf880",
   303 => x"8011740c",
   304 => x"8480808a",
   305 => x"8e04708f",
   306 => x"ffff2491",
   307 => x"3880720c",
   308 => x"8fffff71",
   309 => x"31730c84",
   310 => x"808089ed",
   311 => x"047093ff",
   312 => x"ff249538",
   313 => x"f0808011",
   314 => x"720c8073",
   315 => x"0c83ffff",
   316 => x"740c8480",
   317 => x"808a8e04",
   318 => x"7097ffff",
   319 => x"24903883",
   320 => x"ffff720c",
   321 => x"80730c97",
   322 => x"ffff7131",
   323 => x"740c0290",
   324 => x"050d0402",
   325 => x"e4050d7a",
   326 => x"8480809b",
   327 => x"fc081070",
   328 => x"8480809b",
   329 => x"fc0c7096",
   330 => x"2a708106",
   331 => x"51575757",
   332 => x"74802e8a",
   333 => x"38758107",
   334 => x"8480809b",
   335 => x"fc0c8480",
   336 => x"809bfc08",
   337 => x"70952a70",
   338 => x"81065156",
   339 => x"5674802e",
   340 => x"8a387581",
   341 => x"32848080",
   342 => x"9bfc0c84",
   343 => x"80809bff",
   344 => x"0b848080",
   345 => x"80f52d55",
   346 => x"81967525",
   347 => x"8b38feea",
   348 => x"15558480",
   349 => x"808ae804",
   350 => x"81158480",
   351 => x"809bf455",
   352 => x"8480809b",
   353 => x"f0548480",
   354 => x"809bec53",
   355 => x"7a525584",
   356 => x"808088dd",
   357 => x"2d748429",
   358 => x"19778480",
   359 => x"809bec08",
   360 => x"29882c8c",
   361 => x"1208058c",
   362 => x"120c7784",
   363 => x"80809bf0",
   364 => x"0829882c",
   365 => x"89cc1208",
   366 => x"0589cc12",
   367 => x"0c778480",
   368 => x"809bf408",
   369 => x"29882c93",
   370 => x"8c120805",
   371 => x"938c120c",
   372 => x"55029c05",
   373 => x"0d0402f0",
   374 => x"050d8480",
   375 => x"809bfc08",
   376 => x"9fffff06",
   377 => x"54828053",
   378 => x"73527651",
   379 => x"8480808a",
   380 => x"932d0290",
   381 => x"050d0402",
   382 => x"e8050d84",
   383 => x"19528195",
   384 => x"5684ec12",
   385 => x"089f2c84",
   386 => x"ec13089f",
   387 => x"2c84ec14",
   388 => x"08327072",
   389 => x"318eac15",
   390 => x"089f2c8e",
   391 => x"ac16089f",
   392 => x"2c8eac17",
   393 => x"08327072",
   394 => x"3197ec18",
   395 => x"089f2c97",
   396 => x"ec19089f",
   397 => x"2c97ec1a",
   398 => x"08327072",
   399 => x"318c1b08",
   400 => x"8329881c",
   401 => x"08100590",
   402 => x"1c081011",
   403 => x"70832c8c",
   404 => x"1e083170",
   405 => x"832b5151",
   406 => x"5153515a",
   407 => x"53515853",
   408 => x"51565170",
   409 => x"80258b38",
   410 => x"74713155",
   411 => x"8480808c",
   412 => x"f5047015",
   413 => x"5589cc12",
   414 => x"08832989",
   415 => x"c8130810",
   416 => x"0589d013",
   417 => x"08101170",
   418 => x"832c89cc",
   419 => x"15083170",
   420 => x"832b5151",
   421 => x"51517080",
   422 => x"258b3873",
   423 => x"71315484",
   424 => x"80808da8",
   425 => x"04701454",
   426 => x"938c1208",
   427 => x"83299388",
   428 => x"13081005",
   429 => x"93901308",
   430 => x"10117083",
   431 => x"2c938c15",
   432 => x"08317083",
   433 => x"2b515151",
   434 => x"51708025",
   435 => x"8b387271",
   436 => x"31538480",
   437 => x"808ddb04",
   438 => x"70135372",
   439 => x"882c7081",
   440 => x"ff067688",
   441 => x"2b87fc80",
   442 => x"80067077",
   443 => x"83fe8006",
   444 => x"07707307",
   445 => x"fc0c5153",
   446 => x"ff188415",
   447 => x"55585153",
   448 => x"758025fd",
   449 => x"fc380298",
   450 => x"050d0402",
   451 => x"e8050d78",
   452 => x"84115356",
   453 => x"81955571",
   454 => x"0884e013",
   455 => x"08057270",
   456 => x"8405540c",
   457 => x"ff155574",
   458 => x"8025ec38",
   459 => x"81557484",
   460 => x"29167070",
   461 => x"70840552",
   462 => x"08701011",
   463 => x"fc140810",
   464 => x"11730810",
   465 => x"1170832c",
   466 => x"74317083",
   467 => x"2b84e018",
   468 => x"70089029",
   469 => x"71083170",
   470 => x"842c7384",
   471 => x"2c05720c",
   472 => x"58585151",
   473 => x"51515481",
   474 => x"18585654",
   475 => x"52819675",
   476 => x"25ffbb38",
   477 => x"0298050d",
   478 => x"0402f405",
   479 => x"0d755181",
   480 => x"97537008",
   481 => x"52818072",
   482 => x"258c38ff",
   483 => x"8012710c",
   484 => x"8480808f",
   485 => x"99048071",
   486 => x"0cff1384",
   487 => x"12525372",
   488 => x"8025df38",
   489 => x"028c050d",
   490 => x"0402ec05",
   491 => x"0d775180",
   492 => x"710c8198",
   493 => x"0b84e012",
   494 => x"5455fc13",
   495 => x"08ff8011",
   496 => x"74085452",
   497 => x"54717125",
   498 => x"8c388180",
   499 => x"14730c84",
   500 => x"80808fe9",
   501 => x"04848072",
   502 => x"258c38fc",
   503 => x"8012730c",
   504 => x"8480808f",
   505 => x"e9048073",
   506 => x"0cff15fc",
   507 => x"14545574",
   508 => x"8024c738",
   509 => x"0294050d",
   510 => x"0402f005",
   511 => x"0d848080",
   512 => x"9bfc0870",
   513 => x"81ff0654",
   514 => x"87ffff06",
   515 => x"89808005",
   516 => x"52765184",
   517 => x"80808a93",
   518 => x"2d029005",
   519 => x"0d0402ec",
   520 => x"050d7753",
   521 => x"80730c80",
   522 => x"0b84e014",
   523 => x"0c841354",
   524 => x"81955573",
   525 => x"08bd29fc",
   526 => x"15080584",
   527 => x"15081186",
   528 => x"2a757084",
   529 => x"05570c53",
   530 => x"ff155574",
   531 => x"8025e438",
   532 => x"0294050d",
   533 => x"0402d805",
   534 => x"0d7b84e0",
   535 => x"110884e4",
   536 => x"12087012",
   537 => x"84e81408",
   538 => x"0584ec14",
   539 => x"08055957",
   540 => x"765b5b58",
   541 => x"82577684",
   542 => x"291884e0",
   543 => x"11700884",
   544 => x"e8130819",
   545 => x"70b42988",
   546 => x"2a730c70",
   547 => x"7e317d5f",
   548 => x"5159811a",
   549 => x"5a5b5553",
   550 => x"81957725",
   551 => x"d93802a8",
   552 => x"050d0402",
   553 => x"dc050d7b",
   554 => x"70537b52",
   555 => x"58848080",
   556 => x"87852d77",
   557 => x"57819759",
   558 => x"8480809b",
   559 => x"fc0880ff",
   560 => x"ff068480",
   561 => x"809bf455",
   562 => x"8480809b",
   563 => x"f0548480",
   564 => x"809bec53",
   565 => x"bfff0551",
   566 => x"84808088",
   567 => x"dd2d8480",
   568 => x"809bfc08",
   569 => x"10708480",
   570 => x"809bfc0c",
   571 => x"70962a70",
   572 => x"81065156",
   573 => x"5674802e",
   574 => x"8a387581",
   575 => x"07848080",
   576 => x"9bfc0c84",
   577 => x"80809bfc",
   578 => x"0870952a",
   579 => x"70810651",
   580 => x"56567480",
   581 => x"2e8a3875",
   582 => x"81328480",
   583 => x"809bfc0c",
   584 => x"8480809b",
   585 => x"fc088f06",
   586 => x"8480809b",
   587 => x"ec087129",
   588 => x"902c84ec",
   589 => x"190c8480",
   590 => x"809bf008",
   591 => x"7129902c",
   592 => x"8eac190c",
   593 => x"8480809b",
   594 => x"f4087129",
   595 => x"902c97ec",
   596 => x"190c55ff",
   597 => x"19841858",
   598 => x"59788025",
   599 => x"feda388c",
   600 => x"18518480",
   601 => x"8090d52d",
   602 => x"89cc1851",
   603 => x"84808090",
   604 => x"d52d938c",
   605 => x"18518480",
   606 => x"8090d52d",
   607 => x"02a4050d",
   608 => x"0402d405",
   609 => x"0d7c7e8c",
   610 => x"11705572",
   611 => x"54841308",
   612 => x"585d5956",
   613 => x"742d89cc",
   614 => x"18705376",
   615 => x"52841708",
   616 => x"565a742d",
   617 => x"938c1870",
   618 => x"53765284",
   619 => x"17085659",
   620 => x"742d8480",
   621 => x"809bfc08",
   622 => x"80ffff06",
   623 => x"8480809b",
   624 => x"f4558480",
   625 => x"809bf054",
   626 => x"8480809b",
   627 => x"ec53bfff",
   628 => x"05518480",
   629 => x"8088dd2d",
   630 => x"8480809b",
   631 => x"fc081070",
   632 => x"8480809b",
   633 => x"fc0c7096",
   634 => x"2a708106",
   635 => x"51565674",
   636 => x"802e8a38",
   637 => x"75810784",
   638 => x"80809bfc",
   639 => x"0c848080",
   640 => x"9bfc0870",
   641 => x"952a7081",
   642 => x"06515656",
   643 => x"74802e8a",
   644 => x"38758132",
   645 => x"8480809b",
   646 => x"fc0c8480",
   647 => x"809bfc08",
   648 => x"708f0671",
   649 => x"10708480",
   650 => x"809bfc0c",
   651 => x"70962a70",
   652 => x"81065153",
   653 => x"58585574",
   654 => x"802e8a38",
   655 => x"75810784",
   656 => x"80809bfc",
   657 => x"0c848080",
   658 => x"9bfc0870",
   659 => x"952a7081",
   660 => x"06515656",
   661 => x"74802e8a",
   662 => x"38758132",
   663 => x"8480809b",
   664 => x"fc0c8480",
   665 => x"809bff0b",
   666 => x"84808080",
   667 => x"f52d5581",
   668 => x"9375258b",
   669 => x"38feed15",
   670 => x"55848080",
   671 => x"94ef0474",
   672 => x"84291884",
   673 => x"80809bec",
   674 => x"08782990",
   675 => x"2c84ec12",
   676 => x"0c848080",
   677 => x"9bf00878",
   678 => x"29902c8e",
   679 => x"ac120c84",
   680 => x"80809bf4",
   681 => x"08782990",
   682 => x"2c97ec12",
   683 => x"0c557a51",
   684 => x"84808090",
   685 => x"d52d7951",
   686 => x"84808090",
   687 => x"d52d7851",
   688 => x"84808090",
   689 => x"d52d02ac",
   690 => x"050d0402",
   691 => x"ec050d84",
   692 => x"80809bfc",
   693 => x"087081ff",
   694 => x"065481ff",
   695 => x"ff0680ff",
   696 => x"ff055277",
   697 => x"51848080",
   698 => x"8a932d84",
   699 => x"80809bfc",
   700 => x"08107084",
   701 => x"80809bfc",
   702 => x"0c70962a",
   703 => x"70810651",
   704 => x"55557380",
   705 => x"2e8a3874",
   706 => x"81078480",
   707 => x"809bfc0c",
   708 => x"8480809b",
   709 => x"fc087095",
   710 => x"2a708106",
   711 => x"51555573",
   712 => x"802e8a38",
   713 => x"74813284",
   714 => x"80809bfc",
   715 => x"0c848080",
   716 => x"9bfc0880",
   717 => x"ff068480",
   718 => x"809bf80c",
   719 => x"0294050d",
   720 => x"0402ec05",
   721 => x"0d841852",
   722 => x"81955589",
   723 => x"cc120888",
   724 => x"2c938c13",
   725 => x"08882c8c",
   726 => x"1408882c",
   727 => x"84ec1508",
   728 => x"05565451",
   729 => x"81ff7425",
   730 => x"843881ff",
   731 => x"548eac12",
   732 => x"08115181",
   733 => x"ff712584",
   734 => x"3881ff51",
   735 => x"97ec1208",
   736 => x"135381ff",
   737 => x"73258438",
   738 => x"81ff5373",
   739 => x"902b7188",
   740 => x"2b077074",
   741 => x"07fc0c51",
   742 => x"ff158413",
   743 => x"53557480",
   744 => x"25ffa838",
   745 => x"0294050d",
   746 => x"0402e805",
   747 => x"0d810b84",
   748 => x"80809bf8",
   749 => x"0c848080",
   750 => x"9a980b84",
   751 => x"80809c80",
   752 => x"53705284",
   753 => x"80809a98",
   754 => x"08545572",
   755 => x"2d81c2e6",
   756 => x"0b848080",
   757 => x"9bfc0cff",
   758 => x"56f80854",
   759 => x"73762e80",
   760 => x"e9387384",
   761 => x"2c537285",
   762 => x"2680d038",
   763 => x"72842984",
   764 => x"80809ab4",
   765 => x"05537208",
   766 => x"04848080",
   767 => x"9a985584",
   768 => x"808098bb",
   769 => x"04848080",
   770 => x"99fc5584",
   771 => x"808098bb",
   772 => x"04848080",
   773 => x"99c45584",
   774 => x"808098bb",
   775 => x"04848080",
   776 => x"99a85584",
   777 => x"808098bb",
   778 => x"04848080",
   779 => x"99e05584",
   780 => x"808098bb",
   781 => x"04848080",
   782 => x"998c5573",
   783 => x"8480809c",
   784 => x"80537552",
   785 => x"75085456",
   786 => x"722d8480",
   787 => x"809c8052",
   788 => x"74518c15",
   789 => x"0853722d",
   790 => x"8480809c",
   791 => x"80527451",
   792 => x"90150853",
   793 => x"722d93c3",
   794 => x"54ff8408",
   795 => x"ff155553",
   796 => x"738025f5",
   797 => x"38848080",
   798 => x"97d90400",
   799 => x"00ffffff",
   800 => x"ff00ffff",
   801 => x"ffff00ff",
   802 => x"ffffff00",
   803 => x"400008a3",
   804 => x"4000081e",
   805 => x"40000981",
   806 => x"400003d0",
   807 => x"40000b41",
   808 => x"400007f9",
   809 => x"0000003f",
   810 => x"400008a3",
   811 => x"4000081e",
   812 => x"40000981",
   813 => x"400003d0",
   814 => x"40000b41",
   815 => x"40000acb",
   816 => x"0000003f",
   817 => x"40000385",
   818 => x"4000081e",
   819 => x"40000355",
   820 => x"400003d0",
   821 => x"400002ef",
   822 => x"400005d6",
   823 => x"0000003f",
   824 => x"40000385",
   825 => x"400007a9",
   826 => x"40000355",
   827 => x"400003d0",
   828 => x"400002ef",
   829 => x"400007f9",
   830 => x"0000003f",
   831 => x"40000385",
   832 => x"40000779",
   833 => x"40000355",
   834 => x"400003d0",
   835 => x"400002ef",
   836 => x"400005d6",
   837 => x"0000003f",
   838 => x"40000385",
   839 => x"4000070b",
   840 => x"40000355",
   841 => x"400003d0",
   842 => x"400005f7",
   843 => x"400005d6",
   844 => x"000000ff",
   845 => x"40000bf9",
   846 => x"40000c05",
   847 => x"40000c11",
   848 => x"40000c1d",
   849 => x"40000c29",
   850 => x"40000c35",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

