-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity WS2812B_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end WS2812B_ROM;

architecture arch of WS2812B_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"84808080",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"40000016",
     7 => x"00000000",
     8 => x"84808096",
     9 => x"ec088480",
    10 => x"8096f008",
    11 => x"84808096",
    12 => x"f4088480",
    13 => x"80809808",
    14 => x"2d848080",
    15 => x"96f40c84",
    16 => x"808096f0",
    17 => x"0c848080",
    18 => x"96ec0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"808096c8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"84808096",
    57 => x"ec708480",
    58 => x"80a3f027",
    59 => x"8e388071",
    60 => x"70840553",
    61 => x"0c848080",
    62 => x"81e50484",
    63 => x"8080808c",
    64 => x"51848080",
    65 => x"95a80402",
    66 => x"f8050d73",
    67 => x"52ff8408",
    68 => x"70882a70",
    69 => x"81065151",
    70 => x"5170802e",
    71 => x"f03871ff",
    72 => x"840c7184",
    73 => x"808096ec",
    74 => x"0c028805",
    75 => x"0d0402f0",
    76 => x"050d7553",
    77 => x"80738480",
    78 => x"8080f52d",
    79 => x"7081ff06",
    80 => x"53535470",
    81 => x"742eb138",
    82 => x"7181ff06",
    83 => x"81145452",
    84 => x"ff840870",
    85 => x"882a7081",
    86 => x"06515151",
    87 => x"70802ef0",
    88 => x"3871ff84",
    89 => x"0c811473",
    90 => x"84808080",
    91 => x"f52d7081",
    92 => x"ff065353",
    93 => x"5470d138",
    94 => x"73848080",
    95 => x"96ec0c02",
    96 => x"90050d04",
    97 => x"02f8050d",
    98 => x"ff840870",
    99 => x"892a7081",
   100 => x"06515252",
   101 => x"70802ef0",
   102 => x"387181ff",
   103 => x"06848080",
   104 => x"96ec0c02",
   105 => x"88050d04",
   106 => x"02c4050d",
   107 => x"0280c005",
   108 => x"84808097",
   109 => x"cc5b5680",
   110 => x"76708405",
   111 => x"5808715e",
   112 => x"5e577c70",
   113 => x"84055e08",
   114 => x"58805b77",
   115 => x"982a7888",
   116 => x"2b595372",
   117 => x"8938765e",
   118 => x"84808085",
   119 => x"e3047b80",
   120 => x"2e81d838",
   121 => x"805c7280",
   122 => x"e42ea138",
   123 => x"7280e426",
   124 => x"8e387280",
   125 => x"e32e80f5",
   126 => x"38848080",
   127 => x"84fb0472",
   128 => x"80f32e80",
   129 => x"d0388480",
   130 => x"8084fb04",
   131 => x"75841771",
   132 => x"087e5c56",
   133 => x"57528755",
   134 => x"739c2a74",
   135 => x"842b5552",
   136 => x"71802e83",
   137 => x"38815989",
   138 => x"72258a38",
   139 => x"b7125284",
   140 => x"808084b8",
   141 => x"04b01252",
   142 => x"78802e89",
   143 => x"38715184",
   144 => x"80808287",
   145 => x"2dff1555",
   146 => x"748025cc",
   147 => x"38805484",
   148 => x"80808594",
   149 => x"04758417",
   150 => x"71087054",
   151 => x"5c575284",
   152 => x"808082ae",
   153 => x"2d7b5484",
   154 => x"80808594",
   155 => x"04758417",
   156 => x"71085557",
   157 => x"52848080",
   158 => x"85cb04a5",
   159 => x"51848080",
   160 => x"82872d72",
   161 => x"51848080",
   162 => x"82872d82",
   163 => x"17578480",
   164 => x"8085d604",
   165 => x"73ff1555",
   166 => x"52807225",
   167 => x"b9387970",
   168 => x"81055b84",
   169 => x"808080f5",
   170 => x"2d705253",
   171 => x"84808082",
   172 => x"872d8117",
   173 => x"57848080",
   174 => x"85940472",
   175 => x"a52e0981",
   176 => x"06893881",
   177 => x"5c848080",
   178 => x"85d60472",
   179 => x"51848080",
   180 => x"82872d81",
   181 => x"1757811b",
   182 => x"5b837b25",
   183 => x"fded3872",
   184 => x"fde0387d",
   185 => x"84808096",
   186 => x"ec0c02bc",
   187 => x"050d0402",
   188 => x"f8050d73",
   189 => x"51bd5280",
   190 => x"710c800b",
   191 => x"81f8120c",
   192 => x"ff128412",
   193 => x"52527180",
   194 => x"25ed3802",
   195 => x"88050d04",
   196 => x"02e8050d",
   197 => x"77841153",
   198 => x"56bb5571",
   199 => x"0881f813",
   200 => x"08057270",
   201 => x"8405540c",
   202 => x"ff155574",
   203 => x"8025ec38",
   204 => x"81557484",
   205 => x"29167070",
   206 => x"70840552",
   207 => x"08701011",
   208 => x"fc140810",
   209 => x"11730810",
   210 => x"1170832c",
   211 => x"74317083",
   212 => x"2b81f818",
   213 => x"70089029",
   214 => x"71083170",
   215 => x"842c7384",
   216 => x"2c05720c",
   217 => x"58585151",
   218 => x"51515481",
   219 => x"18585654",
   220 => x"52bc7525",
   221 => x"ffbc3802",
   222 => x"98050d04",
   223 => x"02f4050d",
   224 => x"7451bd53",
   225 => x"70085281",
   226 => x"8072258c",
   227 => x"38ff8012",
   228 => x"710c8480",
   229 => x"80879b04",
   230 => x"80710cff",
   231 => x"13841252",
   232 => x"53728025",
   233 => x"df38028c",
   234 => x"050d0402",
   235 => x"ec050d76",
   236 => x"5180710c",
   237 => x"be0b81f8",
   238 => x"125455fc",
   239 => x"1308ff80",
   240 => x"11740854",
   241 => x"52547171",
   242 => x"258c3881",
   243 => x"8014730c",
   244 => x"84808087",
   245 => x"ea048480",
   246 => x"72258c38",
   247 => x"fc801273",
   248 => x"0c848080",
   249 => x"87ea0480",
   250 => x"730cff15",
   251 => x"fc145455",
   252 => x"748024c7",
   253 => x"38029405",
   254 => x"0d0402ec",
   255 => x"050d7653",
   256 => x"80730c80",
   257 => x"0b81f814",
   258 => x"0c841354",
   259 => x"bb557308",
   260 => x"bd29fc15",
   261 => x"08058415",
   262 => x"0811862a",
   263 => x"75708405",
   264 => x"570c53ff",
   265 => x"15557480",
   266 => x"25e43802",
   267 => x"94050d04",
   268 => x"02f0050d",
   269 => x"7577797b",
   270 => x"57555351",
   271 => x"97ffff71",
   272 => x"258b3870",
   273 => x"1011ffb8",
   274 => x"80801151",
   275 => x"517083ff",
   276 => x"ff248f38",
   277 => x"83ffff72",
   278 => x"0c70730c",
   279 => x"84808088",
   280 => x"f5047087",
   281 => x"ffff2496",
   282 => x"3887ffff",
   283 => x"7131720c",
   284 => x"83ffff73",
   285 => x"0c80740c",
   286 => x"84808089",
   287 => x"e104708b",
   288 => x"ffff2495",
   289 => x"3880720c",
   290 => x"83ffff73",
   291 => x"0cf88080",
   292 => x"11740c84",
   293 => x"808089e1",
   294 => x"04708fff",
   295 => x"ff249138",
   296 => x"80720c8f",
   297 => x"ffff7131",
   298 => x"730c8480",
   299 => x"8089c004",
   300 => x"7093ffff",
   301 => x"249538f0",
   302 => x"80801172",
   303 => x"0c80730c",
   304 => x"83ffff74",
   305 => x"0c848080",
   306 => x"89e10470",
   307 => x"97ffff24",
   308 => x"903883ff",
   309 => x"ff720c80",
   310 => x"730c97ff",
   311 => x"ff713174",
   312 => x"0c029005",
   313 => x"0d0402e4",
   314 => x"050d7984",
   315 => x"80809ffc",
   316 => x"08107084",
   317 => x"80809ffc",
   318 => x"0c70962a",
   319 => x"70810651",
   320 => x"57575774",
   321 => x"802e8a38",
   322 => x"75810784",
   323 => x"80809ffc",
   324 => x"0c848080",
   325 => x"9ffc0870",
   326 => x"952a7081",
   327 => x"06515656",
   328 => x"74802e8a",
   329 => x"38758132",
   330 => x"8480809f",
   331 => x"fc0c8480",
   332 => x"809ffc08",
   333 => x"bf068105",
   334 => x"55bb7525",
   335 => x"8338bb55",
   336 => x"84808098",
   337 => x"94548480",
   338 => x"80989053",
   339 => x"84808098",
   340 => x"8c527851",
   341 => x"84808088",
   342 => x"b02d7482",
   343 => x"2b778480",
   344 => x"80988c08",
   345 => x"29882c84",
   346 => x"8080989c",
   347 => x"12080584",
   348 => x"8080989c",
   349 => x"120c7784",
   350 => x"80809890",
   351 => x"0829882c",
   352 => x"8480809c",
   353 => x"8c120805",
   354 => x"8480809c",
   355 => x"8c120c77",
   356 => x"84808098",
   357 => x"94082988",
   358 => x"2c848080",
   359 => x"a0801208",
   360 => x"05848080",
   361 => x"a080120c",
   362 => x"55029c05",
   363 => x"0d0402f4",
   364 => x"050d8480",
   365 => x"809ffc08",
   366 => x"9fffff06",
   367 => x"53828052",
   368 => x"72518480",
   369 => x"8089e62d",
   370 => x"028c050d",
   371 => x"0402c805",
   372 => x"0d848080",
   373 => x"98980852",
   374 => x"71802e8f",
   375 => x"38ff1284",
   376 => x"80809898",
   377 => x"0c848080",
   378 => x"8c830484",
   379 => x"80808bae",
   380 => x"2d848080",
   381 => x"9fff0b84",
   382 => x"808080f5",
   383 => x"2d848080",
   384 => x"98980c84",
   385 => x"8080a080",
   386 => x"0b840584",
   387 => x"80809c8c",
   388 => x"0b840584",
   389 => x"8080989c",
   390 => x"0b840581",
   391 => x"f81381f8",
   392 => x"1381f813",
   393 => x"5d5d5d5d",
   394 => x"5d5dbb5e",
   395 => x"77089f2c",
   396 => x"78089f2c",
   397 => x"79083270",
   398 => x"72317b08",
   399 => x"9f2c7c08",
   400 => x"9f2c7d08",
   401 => x"32707231",
   402 => x"7f089f2c",
   403 => x"60089f2c",
   404 => x"61083270",
   405 => x"72316370",
   406 => x"70840552",
   407 => x"08701011",
   408 => x"66fc0508",
   409 => x"10117308",
   410 => x"10117083",
   411 => x"2c743170",
   412 => x"832b5151",
   413 => x"5151555e",
   414 => x"5c515c53",
   415 => x"515a5351",
   416 => x"58527180",
   417 => x"258b3876",
   418 => x"72315784",
   419 => x"80808d94",
   420 => x"04711757",
   421 => x"7b707084",
   422 => x"05520870",
   423 => x"1011fc1f",
   424 => x"08101173",
   425 => x"08101170",
   426 => x"832c7431",
   427 => x"70832b56",
   428 => x"51515155",
   429 => x"55527180",
   430 => x"258b3875",
   431 => x"72315684",
   432 => x"80808dc8",
   433 => x"04711656",
   434 => x"7c707084",
   435 => x"05520870",
   436 => x"10117ffc",
   437 => x"05081011",
   438 => x"73081011",
   439 => x"70832c74",
   440 => x"3170832b",
   441 => x"56515151",
   442 => x"55555271",
   443 => x"80258b38",
   444 => x"74723155",
   445 => x"8480808d",
   446 => x"fd047115",
   447 => x"5574882c",
   448 => x"7081ff06",
   449 => x"78882b87",
   450 => x"fc808006",
   451 => x"707983fe",
   452 => x"80060770",
   453 => x"7307fc0c",
   454 => x"51547fff",
   455 => x"05841b84",
   456 => x"1d841f60",
   457 => x"84056284",
   458 => x"05648405",
   459 => x"4543415f",
   460 => x"5d5b4051",
   461 => x"557d8025",
   462 => x"fdf23884",
   463 => x"8080989c",
   464 => x"51848080",
   465 => x"86902d84",
   466 => x"80809c8c",
   467 => x"51848080",
   468 => x"86902d84",
   469 => x"8080a080",
   470 => x"51848080",
   471 => x"86902d02",
   472 => x"b8050d04",
   473 => x"02e4050d",
   474 => x"787a7c57",
   475 => x"57578154",
   476 => x"73822b84",
   477 => x"80809c8c",
   478 => x"1108882c",
   479 => x"848080a0",
   480 => x"80120888",
   481 => x"2c848080",
   482 => x"989c1308",
   483 => x"882c1a53",
   484 => x"55535181",
   485 => x"ff712584",
   486 => x"3881ff51",
   487 => x"75125281",
   488 => x"ff722584",
   489 => x"3881ff52",
   490 => x"74135381",
   491 => x"ff732584",
   492 => x"3881ff53",
   493 => x"70902b72",
   494 => x"882b0770",
   495 => x"7407fc0c",
   496 => x"51811454",
   497 => x"bc7425ff",
   498 => x"a738029c",
   499 => x"050d0402",
   500 => x"f0050d84",
   501 => x"80809898",
   502 => x"08547380",
   503 => x"2e8f38ff",
   504 => x"14848080",
   505 => x"98980c84",
   506 => x"80809081",
   507 => x"04848080",
   508 => x"8bae2d84",
   509 => x"80809ffc",
   510 => x"08bf0684",
   511 => x"80809898",
   512 => x"0c805380",
   513 => x"52805184",
   514 => x"80808ee4",
   515 => x"2d848080",
   516 => x"989c5184",
   517 => x"808086fc",
   518 => x"2d848080",
   519 => x"9c8c5184",
   520 => x"808086fc",
   521 => x"2d848080",
   522 => x"a0805184",
   523 => x"808086fc",
   524 => x"2d029005",
   525 => x"0d0402f0",
   526 => x"050d8480",
   527 => x"80989808",
   528 => x"5473802e",
   529 => x"8f38ff14",
   530 => x"84808098",
   531 => x"980c8480",
   532 => x"8090ec04",
   533 => x"8480808b",
   534 => x"ae2d8480",
   535 => x"809fff0b",
   536 => x"84808080",
   537 => x"f52d8480",
   538 => x"8098980c",
   539 => x"80538052",
   540 => x"80518480",
   541 => x"808ee42d",
   542 => x"84808098",
   543 => x"9c518480",
   544 => x"8087fa2d",
   545 => x"8480809c",
   546 => x"8c518480",
   547 => x"8087fa2d",
   548 => x"848080a0",
   549 => x"80518480",
   550 => x"8087fa2d",
   551 => x"0290050d",
   552 => x"0402ec05",
   553 => x"0d848080",
   554 => x"98980854",
   555 => x"73802e8f",
   556 => x"38ff1484",
   557 => x"80809898",
   558 => x"0c848080",
   559 => x"92a90484",
   560 => x"80809ffc",
   561 => x"087081ff",
   562 => x"06538fff",
   563 => x"ff068880",
   564 => x"80075184",
   565 => x"808089e6",
   566 => x"2d848080",
   567 => x"9ffc0810",
   568 => x"70848080",
   569 => x"9ffc0c70",
   570 => x"962a7081",
   571 => x"06515555",
   572 => x"73802e8a",
   573 => x"38748107",
   574 => x"8480809f",
   575 => x"fc0c8480",
   576 => x"809ffc08",
   577 => x"70952a70",
   578 => x"81065155",
   579 => x"5573802e",
   580 => x"8a387481",
   581 => x"32848080",
   582 => x"9ffc0c84",
   583 => x"80809ffc",
   584 => x"08bf0684",
   585 => x"80809898",
   586 => x"0c805380",
   587 => x"52805184",
   588 => x"80808ee4",
   589 => x"2d848080",
   590 => x"989c5184",
   591 => x"808087ab",
   592 => x"2d848080",
   593 => x"9c8c5184",
   594 => x"808087ab",
   595 => x"2d848080",
   596 => x"a0805184",
   597 => x"808087ab",
   598 => x"2d029405",
   599 => x"0d0402e8",
   600 => x"050d8480",
   601 => x"80989808",
   602 => x"5574802e",
   603 => x"8f38ff15",
   604 => x"84808098",
   605 => x"980c8480",
   606 => x"8093e704",
   607 => x"8480809f",
   608 => x"fc087081",
   609 => x"ff065381",
   610 => x"ffff0680",
   611 => x"ffff0551",
   612 => x"84808089",
   613 => x"e62d8480",
   614 => x"809ffc08",
   615 => x"10708480",
   616 => x"809ffc0c",
   617 => x"70962a70",
   618 => x"81065156",
   619 => x"5674802e",
   620 => x"8a387581",
   621 => x"07848080",
   622 => x"9ffc0c84",
   623 => x"80809ffc",
   624 => x"0870952a",
   625 => x"70810651",
   626 => x"56567480",
   627 => x"2e8a3875",
   628 => x"81328480",
   629 => x"809ffc0c",
   630 => x"8480809f",
   631 => x"fc0880ff",
   632 => x"06848080",
   633 => x"98980c84",
   634 => x"80809ffc",
   635 => x"0880ffff",
   636 => x"06848080",
   637 => x"98945584",
   638 => x"80809890",
   639 => x"54848080",
   640 => x"988c53bf",
   641 => x"ff055184",
   642 => x"808088b0",
   643 => x"2d848080",
   644 => x"9ffc0810",
   645 => x"70848080",
   646 => x"9ffc0c70",
   647 => x"962a7081",
   648 => x"06515656",
   649 => x"74802e8a",
   650 => x"38758107",
   651 => x"8480809f",
   652 => x"fc0c8480",
   653 => x"809ffc08",
   654 => x"70952a70",
   655 => x"81065156",
   656 => x"5674802e",
   657 => x"8a387581",
   658 => x"32848080",
   659 => x"9ffc0c84",
   660 => x"80809ffc",
   661 => x"08830684",
   662 => x"80809894",
   663 => x"08712990",
   664 => x"2c548480",
   665 => x"80989008",
   666 => x"7129902c",
   667 => x"53848080",
   668 => x"988c0871",
   669 => x"29902c52",
   670 => x"55848080",
   671 => x"8ee42d84",
   672 => x"8080989c",
   673 => x"51848080",
   674 => x"87fa2d84",
   675 => x"80809c8c",
   676 => x"51848080",
   677 => x"87fa2d84",
   678 => x"8080a080",
   679 => x"51848080",
   680 => x"87fa2d02",
   681 => x"98050d04",
   682 => x"02f4050d",
   683 => x"810b8480",
   684 => x"8098980c",
   685 => x"84808098",
   686 => x"9c518480",
   687 => x"8085ef2d",
   688 => x"8480809c",
   689 => x"8c518480",
   690 => x"8085ef2d",
   691 => x"848080a0",
   692 => x"80518480",
   693 => x"8085ef2d",
   694 => x"81c2e60b",
   695 => x"8480809f",
   696 => x"fc0cf808",
   697 => x"70842c51",
   698 => x"52718426",
   699 => x"80c43871",
   700 => x"84298480",
   701 => x"8096d805",
   702 => x"52710804",
   703 => x"8480808b",
   704 => x"cd2d8480",
   705 => x"8096b204",
   706 => x"8480808f",
   707 => x"cf2d8480",
   708 => x"8096b204",
   709 => x"84808090",
   710 => x"b62d8480",
   711 => x"8096b204",
   712 => x"84808092",
   713 => x"de2d8480",
   714 => x"8096b204",
   715 => x"84808091",
   716 => x"a12dbacb",
   717 => x"53ff8408",
   718 => x"ff145452",
   719 => x"728025f5",
   720 => x"38848080",
   721 => x"95e20400",
   722 => x"00ffffff",
   723 => x"ff00ffff",
   724 => x"ffff00ff",
   725 => x"ffffff00",
   726 => x"40000afc",
   727 => x"40000b08",
   728 => x"40000b14",
   729 => x"40000b20",
   730 => x"40000b2c",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

