-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity WS2812B_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end WS2812B_ROM;

architecture arch of WS2812B_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"84808080",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"40000016",
     7 => x"00000000",
     8 => x"84808096",
     9 => x"9c088480",
    10 => x"8096a008",
    11 => x"84808096",
    12 => x"a4088480",
    13 => x"80809808",
    14 => x"2d848080",
    15 => x"96a40c84",
    16 => x"808096a0",
    17 => x"0c848080",
    18 => x"969c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"808095f8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"84808096",
    57 => x"9c708480",
    58 => x"80a3a027",
    59 => x"8e388071",
    60 => x"70840553",
    61 => x"0c848080",
    62 => x"81e50484",
    63 => x"8080808c",
    64 => x"51848080",
    65 => x"94d60402",
    66 => x"f8050d73",
    67 => x"52ff8408",
    68 => x"70882a70",
    69 => x"81065151",
    70 => x"5170802e",
    71 => x"f03871ff",
    72 => x"840c7184",
    73 => x"8080969c",
    74 => x"0c028805",
    75 => x"0d0402f0",
    76 => x"050d7553",
    77 => x"80738480",
    78 => x"8080f52d",
    79 => x"7081ff06",
    80 => x"53535470",
    81 => x"742eb138",
    82 => x"7181ff06",
    83 => x"81145452",
    84 => x"ff840870",
    85 => x"882a7081",
    86 => x"06515151",
    87 => x"70802ef0",
    88 => x"3871ff84",
    89 => x"0c811473",
    90 => x"84808080",
    91 => x"f52d7081",
    92 => x"ff065353",
    93 => x"5470d138",
    94 => x"73848080",
    95 => x"969c0c02",
    96 => x"90050d04",
    97 => x"02f8050d",
    98 => x"ff840870",
    99 => x"892a7081",
   100 => x"06515252",
   101 => x"70802ef0",
   102 => x"387181ff",
   103 => x"06848080",
   104 => x"969c0c02",
   105 => x"88050d04",
   106 => x"02c4050d",
   107 => x"0280c005",
   108 => x"84808096",
   109 => x"fc5b5680",
   110 => x"76708405",
   111 => x"5808715e",
   112 => x"5e577c70",
   113 => x"84055e08",
   114 => x"58805b77",
   115 => x"982a7888",
   116 => x"2b595372",
   117 => x"8938765e",
   118 => x"84808085",
   119 => x"e3047b80",
   120 => x"2e81d838",
   121 => x"805c7280",
   122 => x"e42ea138",
   123 => x"7280e426",
   124 => x"8e387280",
   125 => x"e32e80f5",
   126 => x"38848080",
   127 => x"84fb0472",
   128 => x"80f32e80",
   129 => x"d0388480",
   130 => x"8084fb04",
   131 => x"75841771",
   132 => x"087e5c56",
   133 => x"57528755",
   134 => x"739c2a74",
   135 => x"842b5552",
   136 => x"71802e83",
   137 => x"38815989",
   138 => x"72258a38",
   139 => x"b7125284",
   140 => x"808084b8",
   141 => x"04b01252",
   142 => x"78802e89",
   143 => x"38715184",
   144 => x"80808287",
   145 => x"2dff1555",
   146 => x"748025cc",
   147 => x"38805484",
   148 => x"80808594",
   149 => x"04758417",
   150 => x"71087054",
   151 => x"5c575284",
   152 => x"808082ae",
   153 => x"2d7b5484",
   154 => x"80808594",
   155 => x"04758417",
   156 => x"71085557",
   157 => x"52848080",
   158 => x"85cb04a5",
   159 => x"51848080",
   160 => x"82872d72",
   161 => x"51848080",
   162 => x"82872d82",
   163 => x"17578480",
   164 => x"8085d604",
   165 => x"73ff1555",
   166 => x"52807225",
   167 => x"b9387970",
   168 => x"81055b84",
   169 => x"808080f5",
   170 => x"2d705253",
   171 => x"84808082",
   172 => x"872d8117",
   173 => x"57848080",
   174 => x"85940472",
   175 => x"a52e0981",
   176 => x"06893881",
   177 => x"5c848080",
   178 => x"85d60472",
   179 => x"51848080",
   180 => x"82872d81",
   181 => x"1757811b",
   182 => x"5b837b25",
   183 => x"fded3872",
   184 => x"fde0387d",
   185 => x"84808096",
   186 => x"9c0c02bc",
   187 => x"050d0402",
   188 => x"f8050d73",
   189 => x"51bd5280",
   190 => x"710c800b",
   191 => x"81f8120c",
   192 => x"ff128412",
   193 => x"52527180",
   194 => x"25ed3802",
   195 => x"88050d04",
   196 => x"02e8050d",
   197 => x"77841153",
   198 => x"56bb5571",
   199 => x"0881f813",
   200 => x"08057270",
   201 => x"8405540c",
   202 => x"ff155574",
   203 => x"8025ec38",
   204 => x"81557484",
   205 => x"29167070",
   206 => x"70840552",
   207 => x"08701011",
   208 => x"fc140810",
   209 => x"11730810",
   210 => x"1170832c",
   211 => x"74317083",
   212 => x"2b81f818",
   213 => x"70089029",
   214 => x"71083170",
   215 => x"842c7384",
   216 => x"2c05720c",
   217 => x"58585151",
   218 => x"51515481",
   219 => x"18585654",
   220 => x"52bc7525",
   221 => x"ffbc3802",
   222 => x"98050d04",
   223 => x"02f4050d",
   224 => x"7451bd53",
   225 => x"70085281",
   226 => x"8072258c",
   227 => x"38ff8012",
   228 => x"710c8480",
   229 => x"80879b04",
   230 => x"80710cff",
   231 => x"13841252",
   232 => x"53728025",
   233 => x"df38028c",
   234 => x"050d0402",
   235 => x"f0050d75",
   236 => x"5180710c",
   237 => x"be0b81f8",
   238 => x"12535471",
   239 => x"08fc1308",
   240 => x"11822c54",
   241 => x"51707325",
   242 => x"8a387272",
   243 => x"0c848080",
   244 => x"87e70482",
   245 => x"8071258c",
   246 => x"38fe8011",
   247 => x"720c8480",
   248 => x"8087e704",
   249 => x"80720cff",
   250 => x"14fc1353",
   251 => x"54738024",
   252 => x"ca380290",
   253 => x"050d0402",
   254 => x"f4050d74",
   255 => x"5180710c",
   256 => x"800b81f8",
   257 => x"120c8411",
   258 => x"52bb5371",
   259 => x"08882972",
   260 => x"08317084",
   261 => x"29fc1408",
   262 => x"05841408",
   263 => x"11852a74",
   264 => x"70840556",
   265 => x"0c5151ff",
   266 => x"13537280",
   267 => x"25dd3802",
   268 => x"8c050d04",
   269 => x"02f0050d",
   270 => x"7577797b",
   271 => x"57555351",
   272 => x"97ffff71",
   273 => x"258b3870",
   274 => x"1011ffb8",
   275 => x"80801151",
   276 => x"517083ff",
   277 => x"ff248f38",
   278 => x"83ffff72",
   279 => x"0c70730c",
   280 => x"84808088",
   281 => x"f9047087",
   282 => x"ffff2496",
   283 => x"3887ffff",
   284 => x"7131720c",
   285 => x"83ffff73",
   286 => x"0c80740c",
   287 => x"84808089",
   288 => x"e504708b",
   289 => x"ffff2495",
   290 => x"3880720c",
   291 => x"83ffff73",
   292 => x"0cf88080",
   293 => x"11740c84",
   294 => x"808089e5",
   295 => x"04708fff",
   296 => x"ff249138",
   297 => x"80720c8f",
   298 => x"ffff7131",
   299 => x"730c8480",
   300 => x"8089c404",
   301 => x"7093ffff",
   302 => x"249538f0",
   303 => x"80801172",
   304 => x"0c80730c",
   305 => x"83ffff74",
   306 => x"0c848080",
   307 => x"89e50470",
   308 => x"97ffff24",
   309 => x"903883ff",
   310 => x"ff720c80",
   311 => x"730c97ff",
   312 => x"ff713174",
   313 => x"0c029005",
   314 => x"0d0402e4",
   315 => x"050d7984",
   316 => x"80809fac",
   317 => x"08107084",
   318 => x"80809fac",
   319 => x"0c70962a",
   320 => x"70810651",
   321 => x"57575774",
   322 => x"802e8a38",
   323 => x"75810784",
   324 => x"80809fac",
   325 => x"0c848080",
   326 => x"9fac0870",
   327 => x"952a7081",
   328 => x"06515656",
   329 => x"74802e8a",
   330 => x"38758132",
   331 => x"8480809f",
   332 => x"ac0c8480",
   333 => x"809fac08",
   334 => x"bf068105",
   335 => x"55bb7525",
   336 => x"8338bb55",
   337 => x"84808097",
   338 => x"c4548480",
   339 => x"8097c053",
   340 => x"84808097",
   341 => x"bc527851",
   342 => x"84808088",
   343 => x"b42d7482",
   344 => x"2b778480",
   345 => x"8097bc08",
   346 => x"29882c84",
   347 => x"808097cc",
   348 => x"12080584",
   349 => x"808097cc",
   350 => x"120c7784",
   351 => x"808097c0",
   352 => x"0829882c",
   353 => x"8480809b",
   354 => x"bc120805",
   355 => x"8480809b",
   356 => x"bc120c77",
   357 => x"84808097",
   358 => x"c4082988",
   359 => x"2c848080",
   360 => x"9fb01208",
   361 => x"05848080",
   362 => x"9fb0120c",
   363 => x"55029c05",
   364 => x"0d0402f4",
   365 => x"050d8480",
   366 => x"809fac08",
   367 => x"9fffff06",
   368 => x"53828052",
   369 => x"72518480",
   370 => x"8089ea2d",
   371 => x"028c050d",
   372 => x"0402c805",
   373 => x"0d848080",
   374 => x"97c80852",
   375 => x"71802e8f",
   376 => x"38ff1284",
   377 => x"808097c8",
   378 => x"0c848080",
   379 => x"8c870484",
   380 => x"80808bb2",
   381 => x"2d848080",
   382 => x"9faf0b84",
   383 => x"808080f5",
   384 => x"2d848080",
   385 => x"97c80c84",
   386 => x"80809fb0",
   387 => x"0b840584",
   388 => x"80809bbc",
   389 => x"0b840584",
   390 => x"808097cc",
   391 => x"0b840581",
   392 => x"f81381f8",
   393 => x"1381f813",
   394 => x"5d5d5d5d",
   395 => x"5d5dbb5e",
   396 => x"77089f2c",
   397 => x"78089f2c",
   398 => x"79083270",
   399 => x"72317b08",
   400 => x"9f2c7c08",
   401 => x"9f2c7d08",
   402 => x"32707231",
   403 => x"7f089f2c",
   404 => x"60089f2c",
   405 => x"61083270",
   406 => x"72316370",
   407 => x"70840552",
   408 => x"08701011",
   409 => x"66fc0508",
   410 => x"10117308",
   411 => x"10117083",
   412 => x"2c743170",
   413 => x"832b5151",
   414 => x"5151555e",
   415 => x"5c515c53",
   416 => x"515a5351",
   417 => x"58527180",
   418 => x"258b3876",
   419 => x"72315784",
   420 => x"80808d98",
   421 => x"04711757",
   422 => x"7b707084",
   423 => x"05520870",
   424 => x"1011fc1f",
   425 => x"08101173",
   426 => x"08101170",
   427 => x"832c7431",
   428 => x"70832b56",
   429 => x"51515155",
   430 => x"55527180",
   431 => x"258b3875",
   432 => x"72315684",
   433 => x"80808dcc",
   434 => x"04711656",
   435 => x"7c707084",
   436 => x"05520870",
   437 => x"10117ffc",
   438 => x"05081011",
   439 => x"73081011",
   440 => x"70832c74",
   441 => x"3170832b",
   442 => x"56515151",
   443 => x"55555271",
   444 => x"80258b38",
   445 => x"74723155",
   446 => x"8480808e",
   447 => x"81047115",
   448 => x"5574882c",
   449 => x"7081ff06",
   450 => x"78882b87",
   451 => x"fc808006",
   452 => x"707983fe",
   453 => x"80060770",
   454 => x"7307fc0c",
   455 => x"51547fff",
   456 => x"05841b84",
   457 => x"1d841f60",
   458 => x"84056284",
   459 => x"05648405",
   460 => x"4543415f",
   461 => x"5d5b4051",
   462 => x"557d8025",
   463 => x"fdf23884",
   464 => x"808097cc",
   465 => x"51848080",
   466 => x"86902d84",
   467 => x"80809bbc",
   468 => x"51848080",
   469 => x"86902d84",
   470 => x"80809fb0",
   471 => x"51848080",
   472 => x"86902d02",
   473 => x"b8050d04",
   474 => x"02e4050d",
   475 => x"787a7c57",
   476 => x"57578154",
   477 => x"73822b84",
   478 => x"80809bbc",
   479 => x"1108882c",
   480 => x"8480809f",
   481 => x"b0120888",
   482 => x"2c848080",
   483 => x"97cc1308",
   484 => x"882c1a53",
   485 => x"55535181",
   486 => x"ff712584",
   487 => x"3881ff51",
   488 => x"75125281",
   489 => x"ff722584",
   490 => x"3881ff52",
   491 => x"74135381",
   492 => x"ff732584",
   493 => x"3881ff53",
   494 => x"70902b72",
   495 => x"882b0770",
   496 => x"7407fc0c",
   497 => x"51811454",
   498 => x"bc7425ff",
   499 => x"a738029c",
   500 => x"050d0402",
   501 => x"f0050d84",
   502 => x"808097c8",
   503 => x"08547380",
   504 => x"2e8f38ff",
   505 => x"14848080",
   506 => x"97c80c84",
   507 => x"80809085",
   508 => x"04848080",
   509 => x"8bb22d84",
   510 => x"80809fac",
   511 => x"08bf0684",
   512 => x"808097c8",
   513 => x"0c805380",
   514 => x"52805184",
   515 => x"80808ee8",
   516 => x"2d848080",
   517 => x"97cc5184",
   518 => x"808086fc",
   519 => x"2d848080",
   520 => x"9bbc5184",
   521 => x"808086fc",
   522 => x"2d848080",
   523 => x"9fb05184",
   524 => x"808086fc",
   525 => x"2d029005",
   526 => x"0d0402f0",
   527 => x"050d8480",
   528 => x"8097c808",
   529 => x"5473802e",
   530 => x"8f38ff14",
   531 => x"84808097",
   532 => x"c80c8480",
   533 => x"8090f004",
   534 => x"8480808b",
   535 => x"b22d8480",
   536 => x"809faf0b",
   537 => x"84808080",
   538 => x"f52d8480",
   539 => x"8097c80c",
   540 => x"80538052",
   541 => x"80518480",
   542 => x"808ee82d",
   543 => x"84808097",
   544 => x"cc518480",
   545 => x"8087f72d",
   546 => x"8480809b",
   547 => x"bc518480",
   548 => x"8087f72d",
   549 => x"8480809f",
   550 => x"b0518480",
   551 => x"8087f72d",
   552 => x"0290050d",
   553 => x"0402f005",
   554 => x"0d848080",
   555 => x"97c80854",
   556 => x"73802e8f",
   557 => x"38ff1484",
   558 => x"808097c8",
   559 => x"0c848080",
   560 => x"91d70484",
   561 => x"80808bb2",
   562 => x"2d848080",
   563 => x"9fac08bf",
   564 => x"06848080",
   565 => x"97c80c80",
   566 => x"53805280",
   567 => x"51848080",
   568 => x"8ee82d84",
   569 => x"808097cc",
   570 => x"51848080",
   571 => x"87ab2d84",
   572 => x"80809bbc",
   573 => x"51848080",
   574 => x"87ab2d84",
   575 => x"80809fb0",
   576 => x"51848080",
   577 => x"87ab2d02",
   578 => x"90050d04",
   579 => x"02e8050d",
   580 => x"84808097",
   581 => x"c8085574",
   582 => x"802e8f38",
   583 => x"ff158480",
   584 => x"8097c80c",
   585 => x"84808093",
   586 => x"95048480",
   587 => x"809fac08",
   588 => x"7081ff06",
   589 => x"5381ffff",
   590 => x"0680ffff",
   591 => x"05518480",
   592 => x"8089ea2d",
   593 => x"8480809f",
   594 => x"ac081070",
   595 => x"8480809f",
   596 => x"ac0c7096",
   597 => x"2a708106",
   598 => x"51565674",
   599 => x"802e8a38",
   600 => x"75810784",
   601 => x"80809fac",
   602 => x"0c848080",
   603 => x"9fac0870",
   604 => x"952a7081",
   605 => x"06515656",
   606 => x"74802e8a",
   607 => x"38758132",
   608 => x"8480809f",
   609 => x"ac0c8480",
   610 => x"809fac08",
   611 => x"80ff0684",
   612 => x"808097c8",
   613 => x"0c848080",
   614 => x"9fac0880",
   615 => x"ffff0684",
   616 => x"808097c4",
   617 => x"55848080",
   618 => x"97c05484",
   619 => x"808097bc",
   620 => x"53bfff05",
   621 => x"51848080",
   622 => x"88b42d84",
   623 => x"80809fac",
   624 => x"08107084",
   625 => x"80809fac",
   626 => x"0c70962a",
   627 => x"70810651",
   628 => x"56567480",
   629 => x"2e8a3875",
   630 => x"81078480",
   631 => x"809fac0c",
   632 => x"8480809f",
   633 => x"ac087095",
   634 => x"2a708106",
   635 => x"51565674",
   636 => x"802e8a38",
   637 => x"75813284",
   638 => x"80809fac",
   639 => x"0c848080",
   640 => x"9fac0887",
   641 => x"06848080",
   642 => x"97c40871",
   643 => x"29902c54",
   644 => x"84808097",
   645 => x"c0087129",
   646 => x"902c5384",
   647 => x"808097bc",
   648 => x"08712990",
   649 => x"2c525584",
   650 => x"80808ee8",
   651 => x"2d848080",
   652 => x"97cc5184",
   653 => x"808087f7",
   654 => x"2d848080",
   655 => x"9bbc5184",
   656 => x"808087f7",
   657 => x"2d848080",
   658 => x"9fb05184",
   659 => x"808087f7",
   660 => x"2d029805",
   661 => x"0d0402f4",
   662 => x"050d810b",
   663 => x"84808097",
   664 => x"c80c8480",
   665 => x"8097cc51",
   666 => x"84808085",
   667 => x"ef2d8480",
   668 => x"809bbc51",
   669 => x"84808085",
   670 => x"ef2d8480",
   671 => x"809fb051",
   672 => x"84808085",
   673 => x"ef2d81c2",
   674 => x"e60b8480",
   675 => x"809fac0c",
   676 => x"f8087084",
   677 => x"2c515271",
   678 => x"842680c4",
   679 => x"38718429",
   680 => x"84808096",
   681 => x"88055271",
   682 => x"08048480",
   683 => x"808bd12d",
   684 => x"84808095",
   685 => x"e0048480",
   686 => x"808fd32d",
   687 => x"84808095",
   688 => x"e0048480",
   689 => x"8090ba2d",
   690 => x"84808095",
   691 => x"e0048480",
   692 => x"80928c2d",
   693 => x"84808095",
   694 => x"e0048480",
   695 => x"8091a52d",
   696 => x"a78753ff",
   697 => x"8408ff14",
   698 => x"54527280",
   699 => x"25f53884",
   700 => x"80809590",
   701 => x"04000000",
   702 => x"00ffffff",
   703 => x"ff00ffff",
   704 => x"ffff00ff",
   705 => x"ffffff00",
   706 => x"40000aaa",
   707 => x"40000ab6",
   708 => x"40000ac2",
   709 => x"40000ace",
   710 => x"40000ada",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

